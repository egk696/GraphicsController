-- FrameBuffer.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FrameBuffer is
	port (
		address       : in    std_logic_vector(19 downto 0) := (others => '0'); --  avalon_sram_slave.address
		byteenable    : in    std_logic_vector(1 downto 0)  := (others => '0'); --                   .byteenable
		read          : in    std_logic                     := '0';             --                   .read
		write         : in    std_logic                     := '0';             --                   .write
		writedata     : in    std_logic_vector(15 downto 0) := (others => '0'); --                   .writedata
		readdata      : out   std_logic_vector(15 downto 0);                    --                   .readdata
		readdatavalid : out   std_logic;                                        --                   .readdatavalid
		clk           : in    std_logic                     := '0';             --                clk.clk
		SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => '0'); -- external_interface.DQ
		SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    --                   .ADDR
		SRAM_LB_N     : out   std_logic;                                        --                   .LB_N
		SRAM_UB_N     : out   std_logic;                                        --                   .UB_N
		SRAM_CE_N     : out   std_logic;                                        --                   .CE_N
		SRAM_OE_N     : out   std_logic;                                        --                   .OE_N
		SRAM_WE_N     : out   std_logic;                                        --                   .WE_N
		reset         : in    std_logic                     := '0'              --              reset.reset
	);
end entity FrameBuffer;

architecture rtl of FrameBuffer is
	component FrameBuffer_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component FrameBuffer_sram_0;

begin

	sram_0 : component FrameBuffer_sram_0
		port map (
			clk           => clk,           --                clk.clk
			reset         => reset,         --              reset.reset
			SRAM_DQ       => SRAM_DQ,       -- external_interface.export
			SRAM_ADDR     => SRAM_ADDR,     --                   .export
			SRAM_LB_N     => SRAM_LB_N,     --                   .export
			SRAM_UB_N     => SRAM_UB_N,     --                   .export
			SRAM_CE_N     => SRAM_CE_N,     --                   .export
			SRAM_OE_N     => SRAM_OE_N,     --                   .export
			SRAM_WE_N     => SRAM_WE_N,     --                   .export
			address       => address,       --  avalon_sram_slave.address
			byteenable    => byteenable,    --                   .byteenable
			read          => read,          --                   .read
			write         => write,         --                   .write
			writedata     => writedata,     --                   .writedata
			readdata      => readdata,      --                   .readdata
			readdatavalid => readdatavalid  --                   .readdatavalid
		);

end architecture rtl; -- of FrameBuffer
