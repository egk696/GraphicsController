----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01/20/2017 04:12:29 AM
-- Design Name: 
-- Module Name: vga_pack
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package system_config_pack is
	--memory
	constant MEM_ADDRESS_BUS_WIDTH : integer := 32;
	constant MEM_DATA_BUS_WIDTH : integer := 32;
	
end package system_config_pack;

